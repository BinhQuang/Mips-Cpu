library verilog;
use verilog.vl_types.all;
entity cpu_pl_tb is
end cpu_pl_tb;
